//Verilog HDL for "shkim", "AMS_VERILOG" "verilog"


module AMS_VERILOG (input x, output y );
assign y= ~x;
endmodule
