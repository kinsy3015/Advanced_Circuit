magic
tech sky130A
timestamp 1731561380
<< checkpaint >>
rect -755 -750 715 734
<< error_p >>
rect 85 -31 86 -18
<< nwell >>
rect -63 14 62 94
<< pwell >>
rect -64 -69 61 -32
<< nmos >>
rect -32 -65 -23 -35
rect 18 -65 27 -35
<< pmos >>
rect -32 20 -23 50
rect 18 20 27 50
<< ndiff >>
rect -55 -38 -32 -35
rect -55 -48 -52 -38
rect -43 -48 -32 -38
rect -55 -53 -32 -48
rect -55 -63 -52 -53
rect -43 -63 -32 -53
rect -55 -65 -32 -63
rect -23 -65 18 -35
rect 27 -37 50 -35
rect 27 -47 38 -37
rect 47 -47 50 -37
rect 27 -53 50 -47
rect 27 -63 38 -53
rect 47 -63 50 -53
rect 27 -65 50 -63
<< pdiff >>
rect -55 48 -32 50
rect -55 38 -52 48
rect -43 38 -32 48
rect -55 33 -32 38
rect -55 23 -52 33
rect -43 23 -32 33
rect -55 20 -32 23
rect -23 45 18 50
rect -23 35 -4 45
rect 5 35 18 45
rect -23 33 18 35
rect -23 23 -4 33
rect 5 23 18 33
rect -23 20 18 23
rect 27 48 50 50
rect 27 38 38 48
rect 47 38 50 48
rect 27 32 50 38
rect 27 22 38 32
rect 47 22 50 32
rect 27 20 50 22
<< ndiffc >>
rect -52 -48 -43 -38
rect -52 -63 -43 -53
rect 38 -47 47 -37
rect 38 -63 47 -53
<< pdiffc >>
rect -52 38 -43 48
rect -52 23 -43 33
rect 38 38 47 48
rect 38 22 47 32
<< psubdiffcont >>
rect -4 35 5 45
rect -4 23 5 33
rect -36 -106 -18 -94
rect 16 -105 34 -93
<< nsubdiffcont >>
rect -58 73 -49 83
rect -40 73 -31 83
rect -58 61 -49 71
<< poly >>
rect -32 50 -23 53
rect 18 50 27 53
rect -32 8 -23 20
rect -75 -3 -23 8
rect -32 -35 -23 -3
rect 18 -20 27 20
rect 18 -29 66 -20
rect 18 -35 27 -29
rect -32 -68 -23 -65
rect 18 -68 27 -65
<< polycont >>
rect -100 -5 -75 12
rect 66 -31 78 -18
<< locali >>
rect -60 83 55 85
rect -60 73 -58 83
rect -49 73 -40 83
rect -31 73 55 83
rect -60 71 55 73
rect -60 61 -58 71
rect -49 61 55 71
rect -60 60 55 61
rect -55 48 -40 60
rect -55 38 -52 48
rect -43 38 -40 48
rect -55 33 -40 38
rect -55 23 -52 33
rect -43 23 -40 33
rect -55 20 -40 23
rect -10 45 10 50
rect -10 35 -4 45
rect 5 35 10 45
rect -10 33 10 35
rect -10 23 -4 33
rect 5 23 10 33
rect -10 5 10 23
rect 35 48 50 60
rect 35 38 38 48
rect 47 38 50 48
rect 35 32 50 38
rect 35 22 38 32
rect 47 22 50 32
rect 35 20 50 22
rect -10 -15 50 5
rect -55 -38 -40 -35
rect -55 -48 -52 -38
rect -43 -48 -40 -38
rect -55 -53 -40 -48
rect -55 -63 -52 -53
rect -43 -63 -40 -53
rect -55 -89 -40 -63
rect 35 -37 50 -15
rect 35 -47 38 -37
rect 47 -47 50 -37
rect 35 -53 50 -47
rect 35 -63 38 -53
rect 47 -63 50 -53
rect 35 -65 50 -63
rect -65 -93 55 -89
rect -65 -94 16 -93
rect -65 -106 -36 -94
rect -18 -105 16 -94
rect 34 -105 55 -93
rect -18 -106 55 -105
rect -65 -110 55 -106
<< labels >>
rlabel polycont -87 3 -87 3 7 A
rlabel locali -2 73 -2 73 1 vcc
rlabel locali -1 -100 -1 -100 5 gnd
rlabel locali 43 -6 43 -6 3 out
rlabel polycont 74 -24 74 -24 3 B
<< end >>
